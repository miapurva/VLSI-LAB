module tcam(W,N);
input [143:0]W;
output [255:0]N;

wire [255:0]d1[3:0];
assign d1[0][255:0] = 256'd120;
assign d1[1][255:0] = 256'd121;
assign d1[2][255:0] = 256'd122;
assign d1[3][255:0] = 256'd123;
wire [255:0]d2[3:0];
assign d2[0][255:0] = 256'd120;
assign d2[1][255:0] = 256'd121;
assign d2[2][255:0] = 256'd122;
assign d2[3][255:0] = 256'd123;
wire [255:0]d3[3:0];
assign d3[0][255:0] = 256'd120;
assign d3[1][255:0] = 256'd121;
assign d3[2][255:0] = 256'd122;
assign d3[3][255:0] = 256'd123;
wire [255:0]d4[3:0];
assign d4[0][255:0] = 256'd120;
assign d4[1][255:0] = 256'd121;
assign d4[2][255:0] = 256'd122;
assign d4[3][255:0] = 256'd123;
wire [255:0]d5[3:0];
assign d5[0][255:0] = 256'd120;
assign d5[1][255:0] = 256'd121;
assign d5[2][255:0] = 256'd122;
assign d5[3][255:0] = 256'd123;
wire [255:0]d6[3:0];
assign d6[0][255:0] = 256'd120;
assign d6[1][255:0] = 256'd121;
assign d6[2][255:0] = 256'd122;
assign d6[3][255:0] = 256'd123;
wire [255:0]d7[3:0];
assign d7[0][255:0] = 256'd120;
assign d7[1][255:0] = 256'd121;
assign d7[2][255:0] = 256'd122;
assign d7[3][255:0] = 256'd123;
wire [255:0]d8[3:0];
assign d8[0][255:0] = 256'd120;
assign d8[1][255:0] = 256'd121;
assign d8[2][255:0] = 256'd122;
assign d8[3][255:0] = 256'd123;
wire [255:0]d9[3:0];
assign d9[0][255:0] = 256'd120;
assign d9[1][255:0] = 256'd121;
assign d9[2][255:0] = 256'd122;
assign d9[3][255:0] = 256'd123;
wire [255:0]d10[3:0];
assign d10[0][255:0] = 256'd120;
assign d10[1][255:0] = 256'd121;
assign d10[2][255:0] = 256'd122;
assign d10[3][255:0] = 256'd123;
wire [255:0]d11[3:0];
assign d11[0][255:0] = 256'd120;
assign d11[1][255:0] = 256'd121;
assign d11[2][255:0] = 256'd122;
assign d11[3][255:0] = 256'd123;
wire [255:0]d12[3:0];
assign d12[0][255:0] = 256'd120;
assign d12[1][255:0] = 256'd121;
assign d12[2][255:0] = 256'd122;
assign d12[3][255:0] = 256'd123;
wire [255:0]d13[3:0];
assign d13[0][255:0] = 256'd120;
assign d13[1][255:0] = 256'd121;
assign d13[2][255:0] = 256'd122;
assign d13[3][255:0] = 256'd123;
wire [255:0]d14[3:0];
assign d14[0][255:0] = 256'd120;
assign d14[1][255:0] = 256'd121;
assign d14[2][255:0] = 256'd122;
assign d14[3][255:0] = 256'd123;
wire [255:0]d15[3:0];
assign d15[0][255:0] = 256'd120;
assign d15[1][255:0] = 256'd121;
assign d15[2][255:0] = 256'd122;
assign d15[3][255:0] = 256'd123;
wire [255:0]d16[3:0];
assign d16[0][255:0] = 256'd120;
assign d16[1][255:0] = 256'd121;
assign d16[2][255:0] = 256'd122;
assign d16[3][255:0] = 256'd123;
wire [255:0]d17[3:0];
assign d17[0][255:0] = 256'd120;
assign d17[1][255:0] = 256'd121;
assign d17[2][255:0] = 256'd122;
assign d17[3][255:0] = 256'd123;
wire [255:0]d18[3:0];
assign d18[0][255:0] = 256'd120;
assign d18[1][255:0] = 256'd121;
assign d18[2][255:0] = 256'd122;
assign d18[3][255:0] = 256'd123;
wire [255:0]d19[3:0];
assign d19[0][255:0] = 256'd120;
assign d19[1][255:0] = 256'd121;
assign d19[2][255:0] = 256'd122;
assign d19[3][255:0] = 256'd123;
wire [255:0]d20[3:0];
assign d20[0][255:0] = 256'd120;
assign d20[1][255:0] = 256'd121;
assign d20[2][255:0] = 256'd122;
assign d20[3][255:0] = 256'd123;
wire [255:0]d21[3:0];
assign d21[0][255:0] = 256'd120;
assign d21[1][255:0] = 256'd121;
assign d21[2][255:0] = 256'd122;
assign d21[3][255:0] = 256'd123;
wire [255:0]d22[3:0];
assign d22[0][255:0] = 256'd120;
assign d22[1][255:0] = 256'd121;
assign d22[2][255:0] = 256'd122;
assign d22[3][255:0] = 256'd123;
wire [255:0]d23[3:0];
assign d23[0][255:0] = 256'd120;
assign d23[1][255:0] = 256'd121;
assign d23[2][255:0] = 256'd122;
assign d23[3][255:0] = 256'd123;
wire [255:0]d24[3:0];
assign d24[0][255:0] = 256'd120;
assign d24[1][255:0] = 256'd121;
assign d24[2][255:0] = 256'd122;
assign d24[3][255:0] = 256'd123;
wire [255:0]d25[3:0];
assign d25[0][255:0] = 256'd120;
assign d25[1][255:0] = 256'd121;
assign d25[2][255:0] = 256'd122;
assign d25[3][255:0] = 256'd123;
wire [255:0]d26[3:0];
assign d26[0][255:0] = 256'd120;
assign d26[1][255:0] = 256'd121;
assign d26[2][255:0] = 256'd122;
assign d26[3][255:0] = 256'd123;
wire [255:0]d27[3:0];
assign d27[0][255:0] = 256'd120;
assign d27[1][255:0] = 256'd121;
assign d27[2][255:0] = 256'd122;
assign d27[3][255:0] = 256'd123;
wire [255:0]d28[3:0];
assign d28[0][255:0] = 256'd120;
assign d28[1][255:0] = 256'd121;
assign d28[2][255:0] = 256'd122;
assign d28[3][255:0] = 256'd123;
wire [255:0]d29[3:0];
assign d29[0][255:0] = 256'd120;
assign d29[1][255:0] = 256'd121;
assign d29[2][255:0] = 256'd122;
assign d29[3][255:0] = 256'd123;
wire [255:0]d30[3:0];
assign d30[0][255:0] = 256'd120;
assign d30[1][255:0] = 256'd121;
assign d30[2][255:0] = 256'd122;
assign d30[3][255:0] = 256'd123;
wire [255:0]d31[3:0];
assign d31[0][255:0] = 256'd120;
assign d31[1][255:0] = 256'd121;
assign d31[2][255:0] = 256'd122;
assign d31[3][255:0] = 256'd123;
wire [255:0]d32[3:0];
assign d32[0][255:0] = 256'd120;
assign d32[1][255:0] = 256'd121;
assign d32[2][255:0] = 256'd122;
assign d32[3][255:0] = 256'd123;
wire [255:0]d33[3:0];
assign d33[0][255:0] = 256'd120;
assign d33[1][255:0] = 256'd121;
assign d33[2][255:0] = 256'd122;
assign d33[3][255:0] = 256'd123;
wire [255:0]d34[3:0];
assign d34[0][255:0] = 256'd120;
assign d34[1][255:0] = 256'd121;
assign d34[2][255:0] = 256'd122;
assign d34[3][255:0] = 256'd123;
wire [255:0]d35[3:0];
assign d35[0][255:0] = 256'd120;
assign d35[1][255:0] = 256'd121;
assign d35[2][255:0] = 256'd122;
assign d35[3][255:0] = 256'd123;
wire [255:0]d36[3:0];
assign d36[0][255:0] = 256'd120;
assign d36[1][255:0] = 256'd121;
assign d36[2][255:0] = 256'd122;
assign d36[3][255:0] = 256'd123;
wire [255:0]d37[3:0];
assign d37[0][255:0] = 256'd120;
assign d37[1][255:0] = 256'd121;
assign d37[2][255:0] = 256'd122;
assign d37[3][255:0] = 256'd123;
wire [255:0]d38[3:0];
assign d38[0][255:0] = 256'd120;
assign d38[1][255:0] = 256'd121;
assign d38[2][255:0] = 256'd122;
assign d38[3][255:0] = 256'd123;
wire [255:0]d39[3:0];
assign d39[0][255:0] = 256'd120;
assign d39[1][255:0] = 256'd121;
assign d39[2][255:0] = 256'd122;
assign d39[3][255:0] = 256'd123;
wire [255:0]d40[3:0];
assign d40[0][255:0] = 256'd120;
assign d40[1][255:0] = 256'd121;
assign d40[2][255:0] = 256'd122;
assign d40[3][255:0] = 256'd123;
wire [255:0]d41[3:0];
assign d41[0][255:0] = 256'd120;
assign d41[1][255:0] = 256'd121;
assign d41[2][255:0] = 256'd122;
assign d41[3][255:0] = 256'd123;
wire [255:0]d42[3:0];
assign d42[0][255:0] = 256'd120;
assign d42[1][255:0] = 256'd121;
assign d42[2][255:0] = 256'd122;
assign d42[3][255:0] = 256'd123;
wire [255:0]d43[3:0];
assign d43[0][255:0] = 256'd120;
assign d43[1][255:0] = 256'd121;
assign d43[2][255:0] = 256'd122;
assign d43[3][255:0] = 256'd123;
wire [255:0]d44[3:0];
assign d44[0][255:0] = 256'd120;
assign d44[1][255:0] = 256'd121;
assign d44[2][255:0] = 256'd122;
assign d44[3][255:0] = 256'd123;
wire [255:0]d45[3:0];
assign d45[0][255:0] = 256'd120;
assign d45[1][255:0] = 256'd121;
assign d45[2][255:0] = 256'd122;
assign d45[3][255:0] = 256'd123;
wire [255:0]d46[3:0];
assign d46[0][255:0] = 256'd120;
assign d46[1][255:0] = 256'd121;
assign d46[2][255:0] = 256'd122;
assign d46[3][255:0] = 256'd123;
wire [255:0]d47[3:0];
assign d47[0][255:0] = 256'd120;
assign d47[1][255:0] = 256'd121;
assign d47[2][255:0] = 256'd122;
assign d47[3][255:0] = 256'd123;
wire [255:0]d48[3:0];
assign d48[0][255:0] = 256'd120;
assign d48[1][255:0] = 256'd121;
assign d48[2][255:0] = 256'd122;
assign d48[3][255:0] = 256'd123;
wire [255:0]d49[3:0];
assign d49[0][255:0] = 256'd120;
assign d49[1][255:0] = 256'd121;
assign d49[2][255:0] = 256'd122;
assign d49[3][255:0] = 256'd123;
wire [255:0]d50[3:0];
assign d50[0][255:0] = 256'd120;
assign d50[1][255:0] = 256'd121;
assign d50[2][255:0] = 256'd122;
assign d50[3][255:0] = 256'd123;
wire [255:0]d51[3:0];
assign d51[0][255:0] = 256'd120;
assign d51[1][255:0] = 256'd121;
assign d51[2][255:0] = 256'd122;
assign d51[3][255:0] = 256'd123;
wire [255:0]d52[3:0];
assign d52[0][255:0] = 256'd120;
assign d52[1][255:0] = 256'd121;
assign d52[2][255:0] = 256'd122;
assign d52[3][255:0] = 256'd123;
wire [255:0]d53[3:0];
assign d53[0][255:0] = 256'd120;
assign d53[1][255:0] = 256'd121;
assign d53[2][255:0] = 256'd122;
assign d53[3][255:0] = 256'd123;
wire [255:0]d54[3:0];
assign d54[0][255:0] = 256'd120;
assign d54[1][255:0] = 256'd121;
assign d54[2][255:0] = 256'd122;
assign d54[3][255:0] = 256'd123;
wire [255:0]d55[3:0];
assign d55[0][255:0] = 256'd120;
assign d55[1][255:0] = 256'd121;
assign d55[2][255:0] = 256'd122;
assign d55[3][255:0] = 256'd123;
wire [255:0]d56[3:0];
assign d56[0][255:0] = 256'd120;
assign d56[1][255:0] = 256'd121;
assign d56[2][255:0] = 256'd122;
assign d56[3][255:0] = 256'd123;
wire [255:0]d57[3:0];
assign d57[0][255:0] = 256'd120;
assign d57[1][255:0] = 256'd121;
assign d57[2][255:0] = 256'd122;
assign d57[3][255:0] = 256'd123;
wire [255:0]d58[3:0];
assign d58[0][255:0] = 256'd120;
assign d58[1][255:0] = 256'd121;
assign d58[2][255:0] = 256'd122;
assign d58[3][255:0] = 256'd123;
wire [255:0]d59[3:0];
assign d59[0][255:0] = 256'd120;
assign d59[1][255:0] = 256'd121;
assign d59[2][255:0] = 256'd122;
assign d59[3][255:0] = 256'd123;
wire [255:0]d60[3:0];
assign d60[0][255:0] = 256'd120;
assign d60[1][255:0] = 256'd121;
assign d60[2][255:0] = 256'd122;
assign d60[3][255:0] = 256'd123;
wire [255:0]d61[3:0];
assign d61[0][255:0] = 256'd120;
assign d61[1][255:0] = 256'd121;
assign d61[2][255:0] = 256'd122;
assign d61[3][255:0] = 256'd123;
wire [255:0]d62[3:0];
assign d62[0][255:0] = 256'd120;
assign d62[1][255:0] = 256'd121;
assign d62[2][255:0] = 256'd122;
assign d62[3][255:0] = 256'd123;
wire [255:0]d63[3:0];
assign d63[0][255:0] = 256'd120;
assign d63[1][255:0] = 256'd121;
assign d63[2][255:0] = 256'd122;
assign d63[3][255:0] = 256'd123;
wire [255:0]d64[3:0];
assign d64[0][255:0] = 256'd120;
assign d64[1][255:0] = 256'd121;
assign d64[2][255:0] = 256'd122;
assign d64[3][255:0] = 256'd123;
wire [255:0]d65[3:0];
assign d65[0][255:0] = 256'd120;
assign d65[1][255:0] = 256'd121;
assign d65[2][255:0] = 256'd122;
assign d65[3][255:0] = 256'd123;
wire [255:0]d66[3:0];
assign d66[0][255:0] = 256'd120;
assign d66[1][255:0] = 256'd121;
assign d66[2][255:0] = 256'd122;
assign d66[3][255:0] = 256'd123;
wire [255:0]d67[3:0];
assign d67[0][255:0] = 256'd120;
assign d67[1][255:0] = 256'd121;
assign d67[2][255:0] = 256'd122;
assign d67[3][255:0] = 256'd123;
wire [255:0]d68[3:0];
assign d68[0][255:0] = 256'd120;
assign d68[1][255:0] = 256'd121;
assign d68[2][255:0] = 256'd122;
assign d68[3][255:0] = 256'd123;
wire [255:0]d69[3:0];
assign d69[0][255:0] = 256'd120;
assign d69[1][255:0] = 256'd121;
assign d69[2][255:0] = 256'd122;
assign d69[3][255:0] = 256'd123;
wire [255:0]d70[3:0];
assign d70[0][255:0] = 256'd120;
assign d70[1][255:0] = 256'd121;
assign d70[2][255:0] = 256'd122;
assign d70[3][255:0] = 256'd123;
wire [255:0]d71[3:0];
assign d71[0][255:0] = 256'd120;
assign d71[1][255:0] = 256'd121;
assign d71[2][255:0] = 256'd122;
assign d71[3][255:0] = 256'd123;
wire [255:0]d72[3:0];
assign d72[0][255:0] = 256'd120;
assign d72[1][255:0] = 256'd121;
assign d72[2][255:0] = 256'd122;
assign d72[3][255:0] = 256'd123;

wire [255:0]out1;
wire [255:0]out2;
wire [255:0]out3;
wire [255:0]out4;
wire [255:0]out5;
wire [255:0]out6;
wire [255:0]out7;
wire [255:0]out8;
wire [255:0]out9;
wire [255:0]out10;
wire [255:0]out11;
wire [255:0]out12;
wire [255:0]out13;
wire [255:0]out14;
wire [255:0]out15;
wire [255:0]out16;
wire [255:0]out17;
wire [255:0]out18;
wire [255:0]out19;
wire [255:0]out20;
wire [255:0]out21;
wire [255:0]out22;
wire [255:0]out23;
wire [255:0]out24;
wire [255:0]out25;
wire [255:0]out26;
wire [255:0]out27;
wire [255:0]out28;
wire [255:0]out29;
wire [255:0]out30;
wire [255:0]out31;
wire [255:0]out32;
wire [255:0]out33;
wire [255:0]out34;
wire [255:0]out35;
wire [255:0]out36;
wire [255:0]out37;
wire [255:0]out38;
wire [255:0]out39;
wire [255:0]out40;
wire [255:0]out41;
wire [255:0]out42;
wire [255:0]out43;
wire [255:0]out44;
wire [255:0]out45;
wire [255:0]out46;
wire [255:0]out47;
wire [255:0]out48;
wire [255:0]out49;
wire [255:0]out50;
wire [255:0]out51;
wire [255:0]out52;
wire [255:0]out53;
wire [255:0]out54;
wire [255:0]out55;
wire [255:0]out56;
wire [255:0]out57;
wire [255:0]out58;
wire [255:0]out59;
wire [255:0]out60;
wire [255:0]out61;
wire [255:0]out62;
wire [255:0]out63;
wire [255:0]out64;
wire [255:0]out65;
wire [255:0]out66;
wire [255:0]out67;
wire [255:0]out68;
wire [255:0]out69;
wire [255:0]out70;
wire [255:0]out71;
wire [255:0]out72;

integer i1;
mux m1(W[1:0],d1[0],d1[1],d1[2],d1[3],out1);
//assign N[255:0] = out1[255:0];
mux m2(W[3:2],d2[0],d2[1],d2[2],d2[3],out2);
mux m3(W[5:4],d3[0],d3[1],d3[2],d3[3],out3);
mux m4(W[7:6],d4[0],d4[1],d4[2],d4[3],out4);
mux m5(W[9:8],d5[0],d5[1],d5[2],d5[3],out5);
mux m6(W[11:10],d6[0],d6[1],d6[2],d6[3],out6);
mux m7(W[13:12],d7[0],d7[1],d7[2],d7[3],out7);
mux m8(W[15:14],d8[0],d8[1],d8[2],d8[3],out8);
mux m9(W[17:16],d9[0],d9[1],d9[2],d9[3],out9);
mux m10(W[19:18],d10[0],d10[1],d10[2],d10[3],out10);
mux m11(W[21:20],d11[0],d11[1],d11[2],d11[3],out11);
mux m12(W[23:22],d12[0],d12[1],d12[2],d12[3],out12);
mux m13(W[25:24],d13[0],d13[1],d13[2],d13[3],out13);
mux m14(W[27:26],d14[0],d14[1],d14[2],d14[3],out14);
mux m15(W[29:28],d15[0],d15[1],d15[2],d15[3],out15);
mux m16(W[31:30],d16[0],d16[1],d16[2],d16[3],out16);
mux m17(W[33:32],d17[0],d17[1],d17[2],d17[3],out17);
mux m18(W[35:34],d18[0],d18[1],d18[2],d18[3],out18);
mux m19(W[37:36],d19[0],d19[1],d19[2],d19[3],out19);
mux m20(W[39:38],d20[0],d20[1],d20[2],d20[3],out20);
mux m21(W[41:40],d21[0],d21[1],d21[2],d21[3],out21);
mux m22(W[43:42],d22[0],d22[1],d22[2],d22[3],out22);
mux m23(W[45:44],d23[0],d23[1],d23[2],d23[3],out23);
mux m24(W[47:46],d24[0],d24[1],d24[2],d24[3],out24);
mux m25(W[49:48],d25[0],d25[1],d25[2],d25[3],out25);
mux m26(W[51:50],d26[0],d26[1],d26[2],d26[3],out26);
mux m27(W[53:52],d27[0],d27[1],d27[2],d27[3],out27);
mux m28(W[55:54],d28[0],d28[1],d28[2],d28[3],out28);
mux m29(W[57:56],d29[0],d29[1],d29[2],d29[3],out29);
mux m30(W[59:58],d30[0],d30[1],d30[2],d30[3],out30);
mux m31(W[61:60],d31[0],d31[1],d31[2],d31[3],out31);
mux m32(W[63:62],d32[0],d32[1],d32[2],d32[3],out32);
mux m33(W[65:64],d33[0],d33[1],d33[2],d33[3],out33);
mux m34(W[67:66],d34[0],d34[1],d34[2],d34[3],out34);
mux m35(W[69:68],d35[0],d35[1],d35[2],d35[3],out35);
mux m36(W[71:70],d36[0],d36[1],d36[2],d36[3],out36);
mux m37(W[73:72],d37[0],d37[1],d37[2],d37[3],out37);
mux m38(W[75:74],d38[0],d38[1],d38[2],d38[3],out38);
mux m39(W[77:76],d39[0],d39[1],d39[2],d39[3],out39);
mux m40(W[79:78],d40[0],d40[1],d40[2],d40[3],out40);
mux m41(W[81:80],d41[0],d41[1],d41[2],d41[3],out41);
mux m42(W[83:82],d42[0],d42[1],d42[2],d42[3],out42);
mux m43(W[85:84],d43[0],d43[1],d43[2],d43[3],out43);
mux m44(W[87:86],d44[0],d44[1],d44[2],d44[3],out44);
mux m45(W[89:88],d45[0],d45[1],d45[2],d45[3],out45);
mux m46(W[91:90],d46[0],d46[1],d46[2],d46[3],out46);
mux m47(W[93:92],d47[0],d47[1],d47[2],d47[3],out47);
mux m48(W[95:94],d48[0],d48[1],d48[2],d48[3],out48);
mux m49(W[97:96],d49[0],d49[1],d49[2],d49[3],out49);
mux m50(W[99:98],d50[0],d50[1],d50[2],d50[3],out50);
mux m51(W[101:100],d51[0],d51[1],d51[2],d51[3],out51);
mux m52(W[103:102],d52[0],d52[1],d52[2],d52[3],out52);
mux m53(W[105:104],d53[0],d53[1],d53[2],d53[3],out53);
mux m54(W[107:106],d54[0],d54[1],d54[2],d54[3],out54);
mux m55(W[109:108],d55[0],d55[1],d55[2],d55[3],out55);
mux m56(W[111:110],d56[0],d56[1],d56[2],d56[3],out56);
mux m57(W[113:112],d57[0],d57[1],d57[2],d57[3],out57);
mux m58(W[115:114],d58[0],d58[1],d58[2],d58[3],out58);
mux m59(W[117:116],d59[0],d59[1],d59[2],d59[3],out59);
mux m60(W[119:118],d60[0],d60[1],d60[2],d60[3],out60);
mux m61(W[121:120],d61[0],d61[1],d61[2],d61[3],out61);
mux m62(W[123:122],d62[0],d62[1],d62[2],d62[3],out62);
mux m63(W[125:124],d63[0],d63[1],d63[2],d63[3],out63);
mux m64(W[127:126],d64[0],d64[1],d64[2],d64[3],out64);
mux m65(W[129:128],d65[0],d65[1],d65[2],d65[3],out65);
mux m66(W[131:130],d66[0],d66[1],d66[2],d66[3],out66);
mux m67(W[133:132],d67[0],d67[1],d67[2],d67[3],out67);
mux m68(W[135:134],d68[0],d68[1],d68[2],d68[3],out68);
mux m69(W[137:136],d69[0],d69[1],d69[2],d69[3],out69);
mux m70(W[139:138],d70[0],d70[1],d70[2],d70[3],out70);
mux m71(W[141:140],d71[0],d71[1],d71[2],d71[3],out71);
mux m72(W[143:142],d72[0],d72[1],d72[2],d72[3],out72);

wire [255:0]and1;
wire [255:0]and2;
assign and1 = out1 & out2 & out3 & out4 & out5 & out6 & out7 & out8 & out9 & out10 &out11 & out12 & out13 & out14 & out15 & out16 & out17 & out18 & out19 & out20 & out21 & out22 & out23 & out24 & out25 & out26 & out27 & out28 & out29 & out30 & out31 & out32 & out33 & out34 & out35 & out36 & out37 & out38 & out39 & out40 & out41 & out42 & out43 & out44 & out45 & out46 & out47 & out48 & out49 & out50 & out51 & out52 & out53 & out54 & out55 & out56 & out57 & out58 & out59 & out60 & out61 & out62 & out63 & out64 & out65 & out66 & out67 & out68 & out69 & out70 & out71 & out72;
wire u;
pe_256 mn(and1,and2,u);

assign N[255:0] = and1[255:0];
endmodule