module cu(out,in,clk);

input clk;
input [31:0]in;
output [31:0]out;

assign out[31:0]=in[31:0];
endmodule

